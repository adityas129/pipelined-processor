module assign_and(
  input wire x,
  input wire y,
  output wire z
);
  assign z = x & y;
endmodule // and_assign
